// Intial Commit